library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity <entity_name> is

	port
	(
		-- Input ports
		<name>	: in  <type>;
		<name>	: in  <type> := <default_value>;

		-- Inout ports
		<name>	: inout <type>;

		-- Output ports
		<name>	: out <type>;
		<name>	: out <type> := <default_value>
	);
end <entity_name>;


architecture <arch_name> of <entity_name> is



begin

	
end <arch_name>;
