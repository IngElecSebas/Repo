library verilog;
use verilog.vl_types.all;
entity DivFreq_vlg_vec_tst is
end DivFreq_vlg_vec_tst;
