library verilog;
use verilog.vl_types.all;
entity Convertidor_vlg_vec_tst is
end Convertidor_vlg_vec_tst;
