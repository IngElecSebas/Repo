library verilog;
use verilog.vl_types.all;
entity DivFreq50_vlg_check_tst is
    port(
        divided_clk     : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DivFreq50_vlg_check_tst;
