library verilog;
use verilog.vl_types.all;
entity DivFreq50_vlg_vec_tst is
end DivFreq50_vlg_vec_tst;
